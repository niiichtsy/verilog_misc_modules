module adder_subtractor (
)
